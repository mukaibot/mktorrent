sample file 1
