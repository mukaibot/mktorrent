sample file 2
